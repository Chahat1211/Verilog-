module andgate(input1, input2, output1);
	assign output1 = input1 & input2;
endmodule;
