module que10(input a, b, c, e, output reg [15:0] d);
always @(*) begin
    case ({e, a, b, c})
        4'b0000: d = 16'b0000000000000001;
        4'b0001: d = 16'b0000000000000010;
        4'b0010: d = 16'b0000000000000100;
        4'b0011: d = 16'b0000000000001000;
        4'b0100: d = 16'b0000000000010000;
        4'b0101: d = 16'b0000000000100000;
        4'b0110: d = 16'b0000000001000000;
        4'b0111: d = 16'b0000000010000000;
        4'b1000: d = 16'b0000000100000000;
        4'b1001: d = 16'b0000001000000000;
        4'b1010: d = 16'b0000010000000000;
        4'b1011: d = 16'b0000100000000000;
        4'b1100: d = 16'b0001000000000000;
        4'b1101: d = 16'b0010000000000000;
        4'b1110: d = 16'b0100000000000000;
        4'b1111: d = 16'b1000000000000000;
        default: d = 16'b0000000000000000; 
    endcase
end
endmodule

