module and_gate(input1, input2, out);
	assign input1 = 1b'0;
	assign input2 = 2b'1;
	assign output = input1 & input2;
endmodule

